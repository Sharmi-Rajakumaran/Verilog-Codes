module bidirectional_buffer();
  
