module siso();
