module 2_4_decoder_tb();

reg [1:0]i_I_tb;
wire [3:0]o_Y_tb;


integer i;

// Instantiation of the decoder RTL design

  a_4_decoder DUT();
