module 4_1_Mux_tb();
  
  
